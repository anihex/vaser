module vaser
// TilesetInfo stores a summary about a tiled tileset
struct TilesetInfo {
	first_gid int
	source    string
}

module vaser

pub struct KeyMap {
pub:
	key   int
	name  string
	shift bool
	ctrl  bool
	alt   bool
}

module vaser

// Entitier defines what each vaöid entity has to offer
interface Entitier {
	update()
	render()
}

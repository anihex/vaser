module vaser
// Image is used to store the texture-id and the dimensions of the loaded image
struct Image {
	id     u32
	width  f32
	height f32
}

module vaser

interface Scener {
	create()
	input(int, int, int, int)
	update()
	render()
}
